class router_rd_driver extends uvm_driver #(read_xtn);

  `uvm_component_utils(router_rd_driver)

  virtual router_if.RDR_MP vif;
  router_rd_agt_config m_cfg;

  extern function new(string name = "router_rd_driver", uvm_component parent);
  extern function void build_phase(uvm_phase phase);
  extern function void connect_phase(uvm_phase phase);
  extern task run_phase(uvm_phase phase);
  extern task send_to_dut(read_xtn xtn);
  extern function void report_phase(uvm_phase phase);

endclass


function router_rd_driver::new(string name = "router_rd_driver", uvm_component parent);
  super.new(name, parent);
endfunction


function void router_rd_driver::build_phase(uvm_phase phase);
  // call super.build_phase
  super.build_phase(phase);

  // get the config object using uvm_config_db
  if(!uvm_config_db #(router_rd_agt_config)::get(this, "","router_rd_agt_config", m_cfg))
    `uvm_fatal("CONFIG", "cannot get() m_cfg from uvm_config_db. Have you set() it?")
endfunction


function void router_rd_driver::connect_phase(uvm_phase phase);
  vif = m_cfg.vif;
endfunction


task router_rd_driver::run_phase(uvm_phase phase);
 /* @(vif.rdr_cb); //1st clock cycle
  vif.rdr_cb.rst <= 0;
  @(vif.rdr_cb); //2nd clock cycle
  vif.rdr_cb.rst <= 1;*/

  forever
	 begin
    		seq_item_port.get_next_item(req);
    	//	`uvm_info("ROUTER_RD_DRIVER", $sformatf("printing from driver \n 		%s", xtn.sprint()), UVM_LOW)

    		send_to_dut(req);
    		seq_item_port.item_done();
  	end
endtask

/*
task router_rd_driver::send_to_dut(read_xtn xtn);
  // Print the transaction
  `uvm_info("ROUTER_RD_DRIVER", $sformatf("printing from driver \n %s", xtn.sprint()), UVM_LOW)

  @(vif.rdr_cb);
 // while(vif.wdr_cb.busy)//0 it come out, 1 infinty loop 
 // @ (vif.wdr_cb); // wait 1 it comes out, 0 it stays until not busy
  wait(vif.rdr_cb.busy==0);
  vif.rdr_cb.pkt_valid <= 1;

	  vif.rdr_cb.data_in <= xtn.header;
  @ (vif.rdr_cb);

  foreach(xtn.payload_data[i])//payload lenght
  begin
	//  while(vif.wdr_cb.busy)
	// @(vif.wdr_cb);
    wait(vif.rdr_cb.busy==0);
    
    vif.rdr_cb.data_in <= xtn.payload_data[i];
    @ (vif.rdr_cb);
  end

  //while(vif.rdr_cb.busy) @ (vif.wdr_cb);
 wait(vif.rdr_cb.busy==0)

  vif.rdr_cb.pkt_valid <= 0;
  vif.rdr_cb.data_in  <= xtn.parity;
  repeat(2) 
	@ (vif.rdr_cb);

  xtn.err = vif.rdr_cb.error;
  m_cfg.drv_data_count++;
  @ (vif.rdr_cb);

endtask*/


task router_rd_driver::send_to_dut(read_xtn xtn);

  begin
  	// Print the transaction
	  `uvm_info("ROUTER_RD_DRIVER", $sformatf("printing from driver \n %s", xtn.sprint()), UVM_LOW)
	@(vif.rdr_cb);
	wait(vif.rdr_cb.v_out)
	repeat(xtn.no_of_cycles)
	 @(vif.rdr_cb);
	vif.rdr_cb.read_enb <= 1'b1;
	wait(vif.rdr_cb.v_out==0)
	 @(vif.rdr_cb);
	vif.rdr_cb.read_enb <= 1'b0;
	m_cfg.drv_data_count++;
repeat(2)
  @(vif.rdr_cb);
	end
endtask
//UVM REPORT_PHASE

function void router_rd_driver::report_phase(uvm_phase phase);
	`uvm_info(get_type_name(), $sformatf("Report: ROUTER read driver sent %0d transaction", m_cfg.drv_data_count),UVM_LOW)
endfunction

